// UVM agent class