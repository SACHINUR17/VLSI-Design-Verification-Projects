// ALU interface code