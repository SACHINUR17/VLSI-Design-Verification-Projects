// UVM sequence class