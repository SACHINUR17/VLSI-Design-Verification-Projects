// UVM scoreboard class