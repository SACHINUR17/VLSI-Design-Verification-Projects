// UVM test class