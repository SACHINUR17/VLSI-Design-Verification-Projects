// UVM monitor class