// UVM environment class