// UVM transaction class