// UVM driver class