`include "ahb_macros.svh"

package ahb_pkg;
  timeunit 1ns;
  timeprecision 1ps;
  
  import uvm_pkg::*;
  import vutils_pkg::*;

  `include "ahb_types.svh"
  `include "ahb_cfg.svh"
  `include "ahb_seq_item.svh"
  `include "ahb_driver.svh"
  `include "ahb_monitor.svh"
  `include "ahb_sequencer.svh"
  `include "ahb_agent.svh"
  `include "ahb_base_seq.svh"
  `include "ahb_mst_rand_seq.svh"
  `include "ahb_slv_resp_seq.svh"

endpackage // ahb_pkg
