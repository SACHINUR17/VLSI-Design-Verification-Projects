// UVM top testbench